module main_sm ();

main_fsm i_main_sm(
.aclk_i              (  ),
.arstn_i             (  ),
.data_pkt_i          (  ),
.valid_pkt_i         (  ),
.ready_pkt_o         (  ),
.addr_req_o          (  ),
.addr_o              (  ),
.addr_ready_i        (  ),
.valid_s_o           (  ),
.transaction_data_o  (  ),
.cache2cpu_ready_i   (  ),
.pre_hit_i           (  ),
.clr_valid_o         (  ),
.wb_hit_i            (  ),
.wb_r_data_i         (  )
);

endmodule